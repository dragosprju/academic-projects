library verilog;
use verilog.vl_types.all;
entity counter8b_test is
end counter8b_test;
