library verilog;
use verilog.vl_types.all;
entity stack_test2 is
end stack_test2;
