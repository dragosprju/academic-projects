library verilog;
use verilog.vl_types.all;
entity mux8b2c_test is
end mux8b2c_test;
