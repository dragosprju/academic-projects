library verilog;
use verilog.vl_types.all;
entity am2940_test_all is
end am2940_test_all;
