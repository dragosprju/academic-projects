library verilog;
use verilog.vl_types.all;
entity am2940_test4 is
end am2940_test4;
