library verilog;
use verilog.vl_types.all;
entity am2910_test is
end am2910_test;
