library verilog;
use verilog.vl_types.all;
entity reg3b_test is
end reg3b_test;
