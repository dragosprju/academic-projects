library verilog;
use verilog.vl_types.all;
entity sprom_test is
end sprom_test;
