library verilog;
use verilog.vl_types.all;
entity stack_test is
end stack_test;
