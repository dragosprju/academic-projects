module instrdec(instr, ccn, zeror, out);
  input[3:0] instr;
  input ccn, zeror;  
  
  output[10:0] out; 
  reg[10:0] out;
  
  always@(instr or ccn or zeror)
  casex({instr, ccn, zeror})
    // plrc, dec, clear, push, pop, respc, selmux[1:0], pln, mapn, vectn
    6'b0000_xx: out = 11'b001_001_11_011;
    6'b0001_1x: out = 11'b000_000_11_011;
    6'b0001_0x: out = 11'b000_100_00_011;
    6'b0010_xx: out = 11'b000_000_00_101;
    6'b0011_1x: out = 11'b000_000_11_011;
    6'b0011_0x: out = 11'b000_000_00_011;
    6'b0100_1x: out = 11'b100_100_11_011;
    6'b0100_0x: out = 11'b100_100_11_011;
    6'b0101_1x: out = 11'b000_100_01_011;
    6'b0101_0x: out = 11'b000_100_00_011;
    6'b0110_1x: out = 11'b000_000_11_011;
    6'b0110_0x: out = 11'b000_000_00_110;
    6'b0111_1x: out = 11'b000_000_01_011;
    6'b0111_0x: out = 11'b000_000_00_011;
    6'b1000_x0: out = 11'b010_000_10_011;
    6'b1000_x1: out = 11'b000_010_11_011;
    6'b1001_x0: out = 11'b010_000_00_011;
    6'b1001_x1: out = 11'b000_000_11_011;
    6'b1010_1x: out = 11'b000_000_11_011;
    6'b1010_0x: out = 11'b000_010_10_011;
    6'b1011_1x: out = 11'b000_000_11_011;
    6'b1011_0x: out = 11'b000_010_00_011;
    6'b1100_xx: out = 11'b100_000_11_011;
    6'b1101_1x: out = 11'b000_000_10_011;
    6'b1101_0x: out = 11'b000_010_11_011;
    6'b1110_xx: out = 11'b000_000_11_011;
    6'b1111_10: out = 11'b010_000_10_011;
    6'b1111_00: out = 11'b010_010_11_011;
    6'b1111_11: out = 11'b000_010_00_011;
    6'b1111_01: out = 11'b000_010_11_011;
  endcase
endmodule
    
  