library verilog;
use verilog.vl_types.all;
entity am2940_test7 is
end am2940_test7;
