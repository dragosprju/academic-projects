library verilog;
use verilog.vl_types.all;
entity reg8b_test is
end reg8b_test;
