library verilog;
use verilog.vl_types.all;
entity mux12bx4 is
    port(
        A               : in     vl_logic_vector(11 downto 0);
        B               : in     vl_logic_vector(11 downto 0);
        C               : in     vl_logic_vector(11 downto 0);
        D               : in     vl_logic_vector(11 downto 0);
        sel             : in     vl_logic_vector(1 downto 0);
        \out\           : out    vl_logic_vector(11 downto 0)
    );
end mux12bx4;
